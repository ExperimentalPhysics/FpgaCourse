`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:      Ushakov M.V. (EvilLord666)
//
// Create Date:   
// Design Name:   
// Module Name:   
// Project Name:  millet_automate_testbench
// Target Device:  
// Tool versions:  
// Description:   testbench on example of Milley automate design
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
////////////////////////////////////////////////////////////////////////////////

module milley_automate_testbench();

reg [1:0] a;
wire [1:0] b;
reg clk;
reg reset;

milley_automate uut(.clk(clk), .reset(reset), .)

endmodule